library verilog;
use verilog.vl_types.all;
entity mma_top_vlg_tst is
end mma_top_vlg_tst;
